library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.types.all;

entity dataentity is
  port (
    init_data : out full_excitation_vec
  );
end dataentity;

architecture behavioral of dataentity is
begin
init_data(intToTimepoint(0))(0)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(0)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(1)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(1)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(2)(0, 0) <= x"0081";
init_data(intToTimepoint(1))(2)(0, 0) <= x"0081";
init_data(intToTimepoint(0))(3)(0, 0) <= x"0309";
init_data(intToTimepoint(1))(3)(0, 0) <= x"0309";
init_data(intToTimepoint(0))(4)(0, 0) <= x"0747";
init_data(intToTimepoint(1))(4)(0, 0) <= x"0747";
init_data(intToTimepoint(0))(5)(0, 0) <= x"0C9E";
init_data(intToTimepoint(1))(5)(0, 0) <= x"0C9E";
init_data(intToTimepoint(0))(6)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(6)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(7)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(7)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(8)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(8)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(9)(0, 0) <= x"00F5";
init_data(intToTimepoint(1))(9)(0, 0) <= x"00F5";
init_data(intToTimepoint(0))(10)(0, 0) <= x"038E";
init_data(intToTimepoint(1))(10)(0, 0) <= x"038E";
init_data(intToTimepoint(0))(11)(0, 0) <= x"0747";
init_data(intToTimepoint(1))(11)(0, 0) <= x"0747";
init_data(intToTimepoint(0))(12)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(12)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(13)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(13)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(14)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(14)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(15)(0, 0) <= x"0004";
init_data(intToTimepoint(1))(15)(0, 0) <= x"0004";
init_data(intToTimepoint(0))(16)(0, 0) <= x"00F5";
init_data(intToTimepoint(1))(16)(0, 0) <= x"00F5";
init_data(intToTimepoint(0))(17)(0, 0) <= x"0309";
init_data(intToTimepoint(1))(17)(0, 0) <= x"0309";
init_data(intToTimepoint(0))(18)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(18)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(19)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(19)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(20)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(20)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(21)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(21)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(22)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(22)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(23)(0, 0) <= x"0081";
init_data(intToTimepoint(1))(23)(0, 0) <= x"0081";
init_data(intToTimepoint(0))(24)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(24)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(25)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(25)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(26)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(26)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(27)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(27)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(28)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(28)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(29)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(29)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(30)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(30)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(31)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(31)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(32)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(32)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(33)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(33)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(34)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(34)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(35)(0, 0) <= x"0000";
init_data(intToTimepoint(1))(35)(0, 0) <= x"0000";
init_data(intToTimepoint(0))(0)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(0)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(1)(0, 1) <= x"0166";
init_data(intToTimepoint(1))(1)(0, 1) <= x"0166";
init_data(intToTimepoint(0))(2)(0, 1) <= x"05BF";
init_data(intToTimepoint(1))(2)(0, 1) <= x"05BF";
init_data(intToTimepoint(0))(3)(0, 1) <= x"0C9E";
init_data(intToTimepoint(1))(3)(0, 1) <= x"0C9E";
init_data(intToTimepoint(0))(4)(0, 1) <= x"1552";
init_data(intToTimepoint(1))(4)(0, 1) <= x"1552";
init_data(intToTimepoint(0))(5)(0, 1) <= x"1F01";
init_data(intToTimepoint(1))(5)(0, 1) <= x"1F01";
init_data(intToTimepoint(0))(6)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(6)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(7)(0, 1) <= x"0190";
init_data(intToTimepoint(1))(7)(0, 1) <= x"0190";
init_data(intToTimepoint(0))(8)(0, 1) <= x"061C";
init_data(intToTimepoint(1))(8)(0, 1) <= x"061C";
init_data(intToTimepoint(0))(9)(0, 1) <= x"0D30";
init_data(intToTimepoint(1))(9)(0, 1) <= x"0D30";
init_data(intToTimepoint(0))(10)(0, 1) <= x"161C";
init_data(intToTimepoint(1))(10)(0, 1) <= x"161C";
init_data(intToTimepoint(0))(11)(0, 1) <= x"2000";
init_data(intToTimepoint(1))(11)(0, 1) <= x"2000";
init_data(intToTimepoint(0))(12)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(12)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(13)(0, 1) <= x"0166";
init_data(intToTimepoint(1))(13)(0, 1) <= x"0166";
init_data(intToTimepoint(0))(14)(0, 1) <= x"05BF";
init_data(intToTimepoint(1))(14)(0, 1) <= x"05BF";
init_data(intToTimepoint(0))(15)(0, 1) <= x"0C9E";
init_data(intToTimepoint(1))(15)(0, 1) <= x"0C9E";
init_data(intToTimepoint(0))(16)(0, 1) <= x"1552";
init_data(intToTimepoint(1))(16)(0, 1) <= x"1552";
init_data(intToTimepoint(0))(17)(0, 1) <= x"1F01";
init_data(intToTimepoint(1))(17)(0, 1) <= x"1F01";
init_data(intToTimepoint(0))(18)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(18)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(19)(0, 1) <= x"00F5";
init_data(intToTimepoint(1))(19)(0, 1) <= x"00F5";
init_data(intToTimepoint(0))(20)(0, 1) <= x"04BC";
init_data(intToTimepoint(1))(20)(0, 1) <= x"04BC";
init_data(intToTimepoint(0))(21)(0, 1) <= x"0AFD";
init_data(intToTimepoint(1))(21)(0, 1) <= x"0AFD";
init_data(intToTimepoint(0))(22)(0, 1) <= x"1310";
init_data(intToTimepoint(1))(22)(0, 1) <= x"1310";
init_data(intToTimepoint(0))(23)(0, 1) <= x"1C23";
init_data(intToTimepoint(1))(23)(0, 1) <= x"1C23";
init_data(intToTimepoint(0))(24)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(24)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(25)(0, 1) <= x"006A";
init_data(intToTimepoint(1))(25)(0, 1) <= x"006A";
init_data(intToTimepoint(0))(26)(0, 1) <= x"034A";
init_data(intToTimepoint(1))(26)(0, 1) <= x"034A";
init_data(intToTimepoint(0))(27)(0, 1) <= x"0890";
init_data(intToTimepoint(1))(27)(0, 1) <= x"0890";
init_data(intToTimepoint(0))(28)(0, 1) <= x"0FA3";
init_data(intToTimepoint(1))(28)(0, 1) <= x"0FA3";
init_data(intToTimepoint(0))(29)(0, 1) <= x"17BD";
init_data(intToTimepoint(1))(29)(0, 1) <= x"17BD";
init_data(intToTimepoint(0))(30)(0, 1) <= x"0000";
init_data(intToTimepoint(1))(30)(0, 1) <= x"0000";
init_data(intToTimepoint(0))(31)(0, 1) <= x"0009";
init_data(intToTimepoint(1))(31)(0, 1) <= x"0009";
init_data(intToTimepoint(0))(32)(0, 1) <= x"01BE";
init_data(intToTimepoint(1))(32)(0, 1) <= x"01BE";
init_data(intToTimepoint(0))(33)(0, 1) <= x"05BF";
init_data(intToTimepoint(1))(33)(0, 1) <= x"05BF";
init_data(intToTimepoint(0))(34)(0, 1) <= x"0B84";
init_data(intToTimepoint(1))(34)(0, 1) <= x"0B84";
init_data(intToTimepoint(0))(35)(0, 1) <= x"1258";
init_data(intToTimepoint(1))(35)(0, 1) <= x"1258";
init_data(intToTimepoint(0))(0)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(0)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(1)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(1)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(2)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(2)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(3)(0, 2) <= x"0004";
init_data(intToTimepoint(1))(3)(0, 2) <= x"0004";
init_data(intToTimepoint(0))(4)(0, 2) <= x"00F5";
init_data(intToTimepoint(1))(4)(0, 2) <= x"00F5";
init_data(intToTimepoint(0))(5)(0, 2) <= x"0309";
init_data(intToTimepoint(1))(5)(0, 2) <= x"0309";
init_data(intToTimepoint(0))(6)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(6)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(7)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(7)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(8)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(8)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(9)(0, 2) <= x"00F5";
init_data(intToTimepoint(1))(9)(0, 2) <= x"00F5";
init_data(intToTimepoint(0))(10)(0, 2) <= x"038E";
init_data(intToTimepoint(1))(10)(0, 2) <= x"038E";
init_data(intToTimepoint(0))(11)(0, 2) <= x"0747";
init_data(intToTimepoint(1))(11)(0, 2) <= x"0747";
init_data(intToTimepoint(0))(12)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(12)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(13)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(13)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(14)(0, 2) <= x"0081";
init_data(intToTimepoint(1))(14)(0, 2) <= x"0081";
init_data(intToTimepoint(0))(15)(0, 2) <= x"0309";
init_data(intToTimepoint(1))(15)(0, 2) <= x"0309";
init_data(intToTimepoint(0))(16)(0, 2) <= x"0747";
init_data(intToTimepoint(1))(16)(0, 2) <= x"0747";
init_data(intToTimepoint(0))(17)(0, 2) <= x"0C9E";
init_data(intToTimepoint(1))(17)(0, 2) <= x"0C9E";
init_data(intToTimepoint(0))(18)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(18)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(19)(0, 2) <= x"0009";
init_data(intToTimepoint(1))(19)(0, 2) <= x"0009";
init_data(intToTimepoint(0))(20)(0, 2) <= x"01BE";
init_data(intToTimepoint(1))(20)(0, 2) <= x"01BE";
init_data(intToTimepoint(0))(21)(0, 2) <= x"05BF";
init_data(intToTimepoint(1))(21)(0, 2) <= x"05BF";
init_data(intToTimepoint(0))(22)(0, 2) <= x"0B84";
init_data(intToTimepoint(1))(22)(0, 2) <= x"0B84";
init_data(intToTimepoint(0))(23)(0, 2) <= x"1258";
init_data(intToTimepoint(1))(23)(0, 2) <= x"1258";
init_data(intToTimepoint(0))(24)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(24)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(25)(0, 2) <= x"006A";
init_data(intToTimepoint(1))(25)(0, 2) <= x"006A";
init_data(intToTimepoint(0))(26)(0, 2) <= x"034A";
init_data(intToTimepoint(1))(26)(0, 2) <= x"034A";
init_data(intToTimepoint(0))(27)(0, 2) <= x"0890";
init_data(intToTimepoint(1))(27)(0, 2) <= x"0890";
init_data(intToTimepoint(0))(28)(0, 2) <= x"0FA3";
init_data(intToTimepoint(1))(28)(0, 2) <= x"0FA3";
init_data(intToTimepoint(0))(29)(0, 2) <= x"17BD";
init_data(intToTimepoint(1))(29)(0, 2) <= x"17BD";
init_data(intToTimepoint(0))(30)(0, 2) <= x"0000";
init_data(intToTimepoint(1))(30)(0, 2) <= x"0000";
init_data(intToTimepoint(0))(31)(0, 2) <= x"00F5";
init_data(intToTimepoint(1))(31)(0, 2) <= x"00F5";
init_data(intToTimepoint(0))(32)(0, 2) <= x"04BC";
init_data(intToTimepoint(1))(32)(0, 2) <= x"04BC";
init_data(intToTimepoint(0))(33)(0, 2) <= x"0AFD";
init_data(intToTimepoint(1))(33)(0, 2) <= x"0AFD";
init_data(intToTimepoint(0))(34)(0, 2) <= x"1310";
init_data(intToTimepoint(1))(34)(0, 2) <= x"1310";
init_data(intToTimepoint(0))(35)(0, 2) <= x"1C23";
init_data(intToTimepoint(1))(35)(0, 2) <= x"1C23";
init_data(intToTimepoint(0))(0)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(0)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(1)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(1)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(2)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(2)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(3)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(3)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(4)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(4)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(5)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(5)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(6)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(6)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(7)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(7)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(8)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(8)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(9)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(9)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(10)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(10)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(11)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(11)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(12)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(12)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(13)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(13)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(14)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(14)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(15)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(15)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(16)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(16)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(17)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(17)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(18)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(18)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(19)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(19)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(20)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(20)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(21)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(21)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(22)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(22)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(23)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(23)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(24)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(24)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(25)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(25)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(26)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(26)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(27)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(27)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(28)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(28)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(29)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(29)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(30)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(30)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(31)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(31)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(32)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(32)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(33)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(33)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(34)(0, 3) <= x"0000";
init_data(intToTimepoint(1))(34)(0, 3) <= x"0000";
init_data(intToTimepoint(0))(35)(0, 3) <= x"0081";
init_data(intToTimepoint(1))(35)(0, 3) <= x"0081";
init_data(intToTimepoint(0))(0)(1, 0) <= x"1258";
init_data(intToTimepoint(1))(0)(1, 0) <= x"1258";
init_data(intToTimepoint(0))(1)(1, 0) <= x"17BD";
init_data(intToTimepoint(1))(1)(1, 0) <= x"17BD";
init_data(intToTimepoint(0))(2)(1, 0) <= x"1C23";
init_data(intToTimepoint(1))(2)(1, 0) <= x"1C23";
init_data(intToTimepoint(0))(3)(1, 0) <= x"1F01";
init_data(intToTimepoint(1))(3)(1, 0) <= x"1F01";
init_data(intToTimepoint(0))(4)(1, 0) <= x"2000";
init_data(intToTimepoint(1))(4)(1, 0) <= x"2000";
init_data(intToTimepoint(0))(5)(1, 0) <= x"1F01";
init_data(intToTimepoint(1))(5)(1, 0) <= x"1F01";
init_data(intToTimepoint(0))(6)(1, 0) <= x"0B84";
init_data(intToTimepoint(1))(6)(1, 0) <= x"0B84";
init_data(intToTimepoint(0))(7)(1, 0) <= x"0FA3";
init_data(intToTimepoint(1))(7)(1, 0) <= x"0FA3";
init_data(intToTimepoint(0))(8)(1, 0) <= x"1310";
init_data(intToTimepoint(1))(8)(1, 0) <= x"1310";
init_data(intToTimepoint(0))(9)(1, 0) <= x"1552";
init_data(intToTimepoint(1))(9)(1, 0) <= x"1552";
init_data(intToTimepoint(0))(10)(1, 0) <= x"161C";
init_data(intToTimepoint(1))(10)(1, 0) <= x"161C";
init_data(intToTimepoint(0))(11)(1, 0) <= x"1552";
init_data(intToTimepoint(1))(11)(1, 0) <= x"1552";
init_data(intToTimepoint(0))(12)(1, 0) <= x"05BF";
init_data(intToTimepoint(1))(12)(1, 0) <= x"05BF";
init_data(intToTimepoint(0))(13)(1, 0) <= x"0890";
init_data(intToTimepoint(1))(13)(1, 0) <= x"0890";
init_data(intToTimepoint(0))(14)(1, 0) <= x"0AFD";
init_data(intToTimepoint(1))(14)(1, 0) <= x"0AFD";
init_data(intToTimepoint(0))(15)(1, 0) <= x"0C9E";
init_data(intToTimepoint(1))(15)(1, 0) <= x"0C9E";
init_data(intToTimepoint(0))(16)(1, 0) <= x"0D30";
init_data(intToTimepoint(1))(16)(1, 0) <= x"0D30";
init_data(intToTimepoint(0))(17)(1, 0) <= x"0C9E";
init_data(intToTimepoint(1))(17)(1, 0) <= x"0C9E";
init_data(intToTimepoint(0))(18)(1, 0) <= x"01BE";
init_data(intToTimepoint(1))(18)(1, 0) <= x"01BE";
init_data(intToTimepoint(0))(19)(1, 0) <= x"034A";
init_data(intToTimepoint(1))(19)(1, 0) <= x"034A";
init_data(intToTimepoint(0))(20)(1, 0) <= x"04BC";
init_data(intToTimepoint(1))(20)(1, 0) <= x"04BC";
init_data(intToTimepoint(0))(21)(1, 0) <= x"05BF";
init_data(intToTimepoint(1))(21)(1, 0) <= x"05BF";
init_data(intToTimepoint(0))(22)(1, 0) <= x"061C";
init_data(intToTimepoint(1))(22)(1, 0) <= x"061C";
init_data(intToTimepoint(0))(23)(1, 0) <= x"05BF";
init_data(intToTimepoint(1))(23)(1, 0) <= x"05BF";
init_data(intToTimepoint(0))(24)(1, 0) <= x"0009";
init_data(intToTimepoint(1))(24)(1, 0) <= x"0009";
init_data(intToTimepoint(0))(25)(1, 0) <= x"006A";
init_data(intToTimepoint(1))(25)(1, 0) <= x"006A";
init_data(intToTimepoint(0))(26)(1, 0) <= x"00F5";
init_data(intToTimepoint(1))(26)(1, 0) <= x"00F5";
init_data(intToTimepoint(0))(27)(1, 0) <= x"0166";
init_data(intToTimepoint(1))(27)(1, 0) <= x"0166";
init_data(intToTimepoint(0))(28)(1, 0) <= x"0190";
init_data(intToTimepoint(1))(28)(1, 0) <= x"0190";
init_data(intToTimepoint(0))(29)(1, 0) <= x"0166";
init_data(intToTimepoint(1))(29)(1, 0) <= x"0166";
init_data(intToTimepoint(0))(30)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(30)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(31)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(31)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(32)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(32)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(33)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(33)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(34)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(34)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(35)(1, 0) <= x"0000";
init_data(intToTimepoint(1))(35)(1, 0) <= x"0000";
init_data(intToTimepoint(0))(0)(1, 1) <= x"28B4";
init_data(intToTimepoint(1))(0)(1, 1) <= x"28B4";
init_data(intToTimepoint(0))(1)(1, 1) <= x"3177";
init_data(intToTimepoint(1))(1)(1, 1) <= x"3177";
init_data(intToTimepoint(0))(2)(1, 1) <= x"386C";
init_data(intToTimepoint(1))(2)(1, 1) <= x"386C";
init_data(intToTimepoint(0))(3)(1, 1) <= x"3CE4";
init_data(intToTimepoint(1))(3)(1, 1) <= x"3CE4";
init_data(intToTimepoint(0))(4)(1, 1) <= x"3E6F";
init_data(intToTimepoint(1))(4)(1, 1) <= x"3E6F";
init_data(intToTimepoint(0))(5)(1, 1) <= x"3CE4";
init_data(intToTimepoint(1))(5)(1, 1) <= x"3CE4";
init_data(intToTimepoint(0))(6)(1, 1) <= x"29E3";
init_data(intToTimepoint(1))(6)(1, 1) <= x"29E3";
init_data(intToTimepoint(0))(7)(1, 1) <= x"32CF";
init_data(intToTimepoint(1))(7)(1, 1) <= x"32CF";
init_data(intToTimepoint(0))(8)(1, 1) <= x"39E3";
init_data(intToTimepoint(1))(8)(1, 1) <= x"39E3";
init_data(intToTimepoint(0))(9)(1, 1) <= x"3E6F";
init_data(intToTimepoint(1))(9)(1, 1) <= x"3E6F";
init_data(intToTimepoint(0))(10)(1, 1) <= x"4000";
init_data(intToTimepoint(1))(10)(1, 1) <= x"4000";
init_data(intToTimepoint(0))(11)(1, 1) <= x"3E6F";
init_data(intToTimepoint(1))(11)(1, 1) <= x"3E6F";
init_data(intToTimepoint(0))(12)(1, 1) <= x"28B4";
init_data(intToTimepoint(1))(12)(1, 1) <= x"28B4";
init_data(intToTimepoint(0))(13)(1, 1) <= x"3177";
init_data(intToTimepoint(1))(13)(1, 1) <= x"3177";
init_data(intToTimepoint(0))(14)(1, 1) <= x"386C";
init_data(intToTimepoint(1))(14)(1, 1) <= x"386C";
init_data(intToTimepoint(0))(15)(1, 1) <= x"3CE4";
init_data(intToTimepoint(1))(15)(1, 1) <= x"3CE4";
init_data(intToTimepoint(0))(16)(1, 1) <= x"3E6F";
init_data(intToTimepoint(1))(16)(1, 1) <= x"3E6F";
init_data(intToTimepoint(0))(17)(1, 1) <= x"3CE4";
init_data(intToTimepoint(1))(17)(1, 1) <= x"3CE4";
init_data(intToTimepoint(0))(18)(1, 1) <= x"2548";
init_data(intToTimepoint(1))(18)(1, 1) <= x"2548";
init_data(intToTimepoint(0))(19)(1, 1) <= x"2D93";
init_data(intToTimepoint(1))(19)(1, 1) <= x"2D93";
init_data(intToTimepoint(0))(20)(1, 1) <= x"342D";
init_data(intToTimepoint(1))(20)(1, 1) <= x"342D";
init_data(intToTimepoint(0))(21)(1, 1) <= x"386C";
init_data(intToTimepoint(1))(21)(1, 1) <= x"386C";
init_data(intToTimepoint(0))(22)(1, 1) <= x"39E3";
init_data(intToTimepoint(1))(22)(1, 1) <= x"39E3";
init_data(intToTimepoint(0))(23)(1, 1) <= x"386C";
init_data(intToTimepoint(1))(23)(1, 1) <= x"386C";
init_data(intToTimepoint(0))(24)(1, 1) <= x"2000";
init_data(intToTimepoint(1))(24)(1, 1) <= x"2000";
init_data(intToTimepoint(0))(25)(1, 1) <= x"278A";
init_data(intToTimepoint(1))(25)(1, 1) <= x"278A";
init_data(intToTimepoint(0))(26)(1, 1) <= x"2D93";
init_data(intToTimepoint(1))(26)(1, 1) <= x"2D93";
init_data(intToTimepoint(0))(27)(1, 1) <= x"3177";
init_data(intToTimepoint(1))(27)(1, 1) <= x"3177";
init_data(intToTimepoint(0))(28)(1, 1) <= x"32CF";
init_data(intToTimepoint(1))(28)(1, 1) <= x"32CF";
init_data(intToTimepoint(0))(29)(1, 1) <= x"3177";
init_data(intToTimepoint(1))(29)(1, 1) <= x"3177";
init_data(intToTimepoint(0))(30)(1, 1) <= x"1971";
init_data(intToTimepoint(1))(30)(1, 1) <= x"1971";
init_data(intToTimepoint(0))(31)(1, 1) <= x"2000";
init_data(intToTimepoint(1))(31)(1, 1) <= x"2000";
init_data(intToTimepoint(0))(32)(1, 1) <= x"2548";
init_data(intToTimepoint(1))(32)(1, 1) <= x"2548";
init_data(intToTimepoint(0))(33)(1, 1) <= x"28B4";
init_data(intToTimepoint(1))(33)(1, 1) <= x"28B4";
init_data(intToTimepoint(0))(34)(1, 1) <= x"29E3";
init_data(intToTimepoint(1))(34)(1, 1) <= x"29E3";
init_data(intToTimepoint(0))(35)(1, 1) <= x"28B4";
init_data(intToTimepoint(1))(35)(1, 1) <= x"28B4";
init_data(intToTimepoint(0))(0)(1, 2) <= x"05BF";
init_data(intToTimepoint(1))(0)(1, 2) <= x"05BF";
init_data(intToTimepoint(0))(1)(1, 2) <= x"0890";
init_data(intToTimepoint(1))(1)(1, 2) <= x"0890";
init_data(intToTimepoint(0))(2)(1, 2) <= x"0AFD";
init_data(intToTimepoint(1))(2)(1, 2) <= x"0AFD";
init_data(intToTimepoint(0))(3)(1, 2) <= x"0C9E";
init_data(intToTimepoint(1))(3)(1, 2) <= x"0C9E";
init_data(intToTimepoint(0))(4)(1, 2) <= x"0D30";
init_data(intToTimepoint(1))(4)(1, 2) <= x"0D30";
init_data(intToTimepoint(0))(5)(1, 2) <= x"0C9E";
init_data(intToTimepoint(1))(5)(1, 2) <= x"0C9E";
init_data(intToTimepoint(0))(6)(1, 2) <= x"0B84";
init_data(intToTimepoint(1))(6)(1, 2) <= x"0B84";
init_data(intToTimepoint(0))(7)(1, 2) <= x"0FA3";
init_data(intToTimepoint(1))(7)(1, 2) <= x"0FA3";
init_data(intToTimepoint(0))(8)(1, 2) <= x"1310";
init_data(intToTimepoint(1))(8)(1, 2) <= x"1310";
init_data(intToTimepoint(0))(9)(1, 2) <= x"1552";
init_data(intToTimepoint(1))(9)(1, 2) <= x"1552";
init_data(intToTimepoint(0))(10)(1, 2) <= x"161C";
init_data(intToTimepoint(1))(10)(1, 2) <= x"161C";
init_data(intToTimepoint(0))(11)(1, 2) <= x"1552";
init_data(intToTimepoint(1))(11)(1, 2) <= x"1552";
init_data(intToTimepoint(0))(12)(1, 2) <= x"1258";
init_data(intToTimepoint(1))(12)(1, 2) <= x"1258";
init_data(intToTimepoint(0))(13)(1, 2) <= x"17BD";
init_data(intToTimepoint(1))(13)(1, 2) <= x"17BD";
init_data(intToTimepoint(0))(14)(1, 2) <= x"1C23";
init_data(intToTimepoint(1))(14)(1, 2) <= x"1C23";
init_data(intToTimepoint(0))(15)(1, 2) <= x"1F01";
init_data(intToTimepoint(1))(15)(1, 2) <= x"1F01";
init_data(intToTimepoint(0))(16)(1, 2) <= x"2000";
init_data(intToTimepoint(1))(16)(1, 2) <= x"2000";
init_data(intToTimepoint(0))(17)(1, 2) <= x"1F01";
init_data(intToTimepoint(1))(17)(1, 2) <= x"1F01";
init_data(intToTimepoint(0))(18)(1, 2) <= x"1971";
init_data(intToTimepoint(1))(18)(1, 2) <= x"1971";
init_data(intToTimepoint(0))(19)(1, 2) <= x"2000";
init_data(intToTimepoint(1))(19)(1, 2) <= x"2000";
init_data(intToTimepoint(0))(20)(1, 2) <= x"2548";
init_data(intToTimepoint(1))(20)(1, 2) <= x"2548";
init_data(intToTimepoint(0))(21)(1, 2) <= x"28B4";
init_data(intToTimepoint(1))(21)(1, 2) <= x"28B4";
init_data(intToTimepoint(0))(22)(1, 2) <= x"29E3";
init_data(intToTimepoint(1))(22)(1, 2) <= x"29E3";
init_data(intToTimepoint(0))(23)(1, 2) <= x"28B4";
init_data(intToTimepoint(1))(23)(1, 2) <= x"28B4";
init_data(intToTimepoint(0))(24)(1, 2) <= x"2000";
init_data(intToTimepoint(1))(24)(1, 2) <= x"2000";
init_data(intToTimepoint(0))(25)(1, 2) <= x"278A";
init_data(intToTimepoint(1))(25)(1, 2) <= x"278A";
init_data(intToTimepoint(0))(26)(1, 2) <= x"2D93";
init_data(intToTimepoint(1))(26)(1, 2) <= x"2D93";
init_data(intToTimepoint(0))(27)(1, 2) <= x"3177";
init_data(intToTimepoint(1))(27)(1, 2) <= x"3177";
init_data(intToTimepoint(0))(28)(1, 2) <= x"32CF";
init_data(intToTimepoint(1))(28)(1, 2) <= x"32CF";
init_data(intToTimepoint(0))(29)(1, 2) <= x"3177";
init_data(intToTimepoint(1))(29)(1, 2) <= x"3177";
init_data(intToTimepoint(0))(30)(1, 2) <= x"2548";
init_data(intToTimepoint(1))(30)(1, 2) <= x"2548";
init_data(intToTimepoint(0))(31)(1, 2) <= x"2D93";
init_data(intToTimepoint(1))(31)(1, 2) <= x"2D93";
init_data(intToTimepoint(0))(32)(1, 2) <= x"342D";
init_data(intToTimepoint(1))(32)(1, 2) <= x"342D";
init_data(intToTimepoint(0))(33)(1, 2) <= x"386C";
init_data(intToTimepoint(1))(33)(1, 2) <= x"386C";
init_data(intToTimepoint(0))(34)(1, 2) <= x"39E3";
init_data(intToTimepoint(1))(34)(1, 2) <= x"39E3";
init_data(intToTimepoint(0))(35)(1, 2) <= x"386C";
init_data(intToTimepoint(1))(35)(1, 2) <= x"386C";
init_data(intToTimepoint(0))(0)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(0)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(1)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(1)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(2)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(2)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(3)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(3)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(4)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(4)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(5)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(5)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(6)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(6)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(7)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(7)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(8)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(8)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(9)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(9)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(10)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(10)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(11)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(11)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(12)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(12)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(13)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(13)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(14)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(14)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(15)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(15)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(16)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(16)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(17)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(17)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(18)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(18)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(19)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(19)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(20)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(20)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(21)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(21)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(22)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(22)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(23)(1, 3) <= x"0000";
init_data(intToTimepoint(1))(23)(1, 3) <= x"0000";
init_data(intToTimepoint(0))(24)(1, 3) <= x"0009";
init_data(intToTimepoint(1))(24)(1, 3) <= x"0009";
init_data(intToTimepoint(0))(25)(1, 3) <= x"006A";
init_data(intToTimepoint(1))(25)(1, 3) <= x"006A";
init_data(intToTimepoint(0))(26)(1, 3) <= x"00F5";
init_data(intToTimepoint(1))(26)(1, 3) <= x"00F5";
init_data(intToTimepoint(0))(27)(1, 3) <= x"0166";
init_data(intToTimepoint(1))(27)(1, 3) <= x"0166";
init_data(intToTimepoint(0))(28)(1, 3) <= x"0190";
init_data(intToTimepoint(1))(28)(1, 3) <= x"0190";
init_data(intToTimepoint(0))(29)(1, 3) <= x"0166";
init_data(intToTimepoint(1))(29)(1, 3) <= x"0166";
init_data(intToTimepoint(0))(30)(1, 3) <= x"01BE";
init_data(intToTimepoint(1))(30)(1, 3) <= x"01BE";
init_data(intToTimepoint(0))(31)(1, 3) <= x"034A";
init_data(intToTimepoint(1))(31)(1, 3) <= x"034A";
init_data(intToTimepoint(0))(32)(1, 3) <= x"04BC";
init_data(intToTimepoint(1))(32)(1, 3) <= x"04BC";
init_data(intToTimepoint(0))(33)(1, 3) <= x"05BF";
init_data(intToTimepoint(1))(33)(1, 3) <= x"05BF";
init_data(intToTimepoint(0))(34)(1, 3) <= x"061C";
init_data(intToTimepoint(1))(34)(1, 3) <= x"061C";
init_data(intToTimepoint(0))(35)(1, 3) <= x"05BF";
init_data(intToTimepoint(1))(35)(1, 3) <= x"05BF";
init_data(intToTimepoint(0))(0)(2, 0) <= x"1C23";
init_data(intToTimepoint(1))(0)(2, 0) <= x"1C23";
init_data(intToTimepoint(0))(1)(2, 0) <= x"17BD";
init_data(intToTimepoint(1))(1)(2, 0) <= x"17BD";
init_data(intToTimepoint(0))(2)(2, 0) <= x"1258";
init_data(intToTimepoint(1))(2)(2, 0) <= x"1258";
init_data(intToTimepoint(0))(3)(2, 0) <= x"0C9E";
init_data(intToTimepoint(1))(3)(2, 0) <= x"0C9E";
init_data(intToTimepoint(0))(4)(2, 0) <= x"0747";
init_data(intToTimepoint(1))(4)(2, 0) <= x"0747";
init_data(intToTimepoint(0))(5)(2, 0) <= x"0309";
init_data(intToTimepoint(1))(5)(2, 0) <= x"0309";
init_data(intToTimepoint(0))(6)(2, 0) <= x"1310";
init_data(intToTimepoint(1))(6)(2, 0) <= x"1310";
init_data(intToTimepoint(0))(7)(2, 0) <= x"0FA3";
init_data(intToTimepoint(1))(7)(2, 0) <= x"0FA3";
init_data(intToTimepoint(0))(8)(2, 0) <= x"0B84";
init_data(intToTimepoint(1))(8)(2, 0) <= x"0B84";
init_data(intToTimepoint(0))(9)(2, 0) <= x"0747";
init_data(intToTimepoint(1))(9)(2, 0) <= x"0747";
init_data(intToTimepoint(0))(10)(2, 0) <= x"038E";
init_data(intToTimepoint(1))(10)(2, 0) <= x"038E";
init_data(intToTimepoint(0))(11)(2, 0) <= x"00F5";
init_data(intToTimepoint(1))(11)(2, 0) <= x"00F5";
init_data(intToTimepoint(0))(12)(2, 0) <= x"0AFD";
init_data(intToTimepoint(1))(12)(2, 0) <= x"0AFD";
init_data(intToTimepoint(0))(13)(2, 0) <= x"0890";
init_data(intToTimepoint(1))(13)(2, 0) <= x"0890";
init_data(intToTimepoint(0))(14)(2, 0) <= x"05BF";
init_data(intToTimepoint(1))(14)(2, 0) <= x"05BF";
init_data(intToTimepoint(0))(15)(2, 0) <= x"0309";
init_data(intToTimepoint(1))(15)(2, 0) <= x"0309";
init_data(intToTimepoint(0))(16)(2, 0) <= x"00F5";
init_data(intToTimepoint(1))(16)(2, 0) <= x"00F5";
init_data(intToTimepoint(0))(17)(2, 0) <= x"0004";
init_data(intToTimepoint(1))(17)(2, 0) <= x"0004";
init_data(intToTimepoint(0))(18)(2, 0) <= x"04BC";
init_data(intToTimepoint(1))(18)(2, 0) <= x"04BC";
init_data(intToTimepoint(0))(19)(2, 0) <= x"034A";
init_data(intToTimepoint(1))(19)(2, 0) <= x"034A";
init_data(intToTimepoint(0))(20)(2, 0) <= x"01BE";
init_data(intToTimepoint(1))(20)(2, 0) <= x"01BE";
init_data(intToTimepoint(0))(21)(2, 0) <= x"0081";
init_data(intToTimepoint(1))(21)(2, 0) <= x"0081";
init_data(intToTimepoint(0))(22)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(22)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(23)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(23)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(24)(2, 0) <= x"00F5";
init_data(intToTimepoint(1))(24)(2, 0) <= x"00F5";
init_data(intToTimepoint(0))(25)(2, 0) <= x"006A";
init_data(intToTimepoint(1))(25)(2, 0) <= x"006A";
init_data(intToTimepoint(0))(26)(2, 0) <= x"0009";
init_data(intToTimepoint(1))(26)(2, 0) <= x"0009";
init_data(intToTimepoint(0))(27)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(27)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(28)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(28)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(29)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(29)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(30)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(30)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(31)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(31)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(32)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(32)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(33)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(33)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(34)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(34)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(35)(2, 0) <= x"0000";
init_data(intToTimepoint(1))(35)(2, 0) <= x"0000";
init_data(intToTimepoint(0))(0)(2, 1) <= x"386C";
init_data(intToTimepoint(1))(0)(2, 1) <= x"386C";
init_data(intToTimepoint(0))(1)(2, 1) <= x"3177";
init_data(intToTimepoint(1))(1)(2, 1) <= x"3177";
init_data(intToTimepoint(0))(2)(2, 1) <= x"28B4";
init_data(intToTimepoint(1))(2)(2, 1) <= x"28B4";
init_data(intToTimepoint(0))(3)(2, 1) <= x"1F01";
init_data(intToTimepoint(1))(3)(2, 1) <= x"1F01";
init_data(intToTimepoint(0))(4)(2, 1) <= x"1552";
init_data(intToTimepoint(1))(4)(2, 1) <= x"1552";
init_data(intToTimepoint(0))(5)(2, 1) <= x"0C9E";
init_data(intToTimepoint(1))(5)(2, 1) <= x"0C9E";
init_data(intToTimepoint(0))(6)(2, 1) <= x"39E3";
init_data(intToTimepoint(1))(6)(2, 1) <= x"39E3";
init_data(intToTimepoint(0))(7)(2, 1) <= x"32CF";
init_data(intToTimepoint(1))(7)(2, 1) <= x"32CF";
init_data(intToTimepoint(0))(8)(2, 1) <= x"29E3";
init_data(intToTimepoint(1))(8)(2, 1) <= x"29E3";
init_data(intToTimepoint(0))(9)(2, 1) <= x"2000";
init_data(intToTimepoint(1))(9)(2, 1) <= x"2000";
init_data(intToTimepoint(0))(10)(2, 1) <= x"161C";
init_data(intToTimepoint(1))(10)(2, 1) <= x"161C";
init_data(intToTimepoint(0))(11)(2, 1) <= x"0D30";
init_data(intToTimepoint(1))(11)(2, 1) <= x"0D30";
init_data(intToTimepoint(0))(12)(2, 1) <= x"386C";
init_data(intToTimepoint(1))(12)(2, 1) <= x"386C";
init_data(intToTimepoint(0))(13)(2, 1) <= x"3177";
init_data(intToTimepoint(1))(13)(2, 1) <= x"3177";
init_data(intToTimepoint(0))(14)(2, 1) <= x"28B4";
init_data(intToTimepoint(1))(14)(2, 1) <= x"28B4";
init_data(intToTimepoint(0))(15)(2, 1) <= x"1F01";
init_data(intToTimepoint(1))(15)(2, 1) <= x"1F01";
init_data(intToTimepoint(0))(16)(2, 1) <= x"1552";
init_data(intToTimepoint(1))(16)(2, 1) <= x"1552";
init_data(intToTimepoint(0))(17)(2, 1) <= x"0C9E";
init_data(intToTimepoint(1))(17)(2, 1) <= x"0C9E";
init_data(intToTimepoint(0))(18)(2, 1) <= x"342D";
init_data(intToTimepoint(1))(18)(2, 1) <= x"342D";
init_data(intToTimepoint(0))(19)(2, 1) <= x"2D93";
init_data(intToTimepoint(1))(19)(2, 1) <= x"2D93";
init_data(intToTimepoint(0))(20)(2, 1) <= x"2548";
init_data(intToTimepoint(1))(20)(2, 1) <= x"2548";
init_data(intToTimepoint(0))(21)(2, 1) <= x"1C23";
init_data(intToTimepoint(1))(21)(2, 1) <= x"1C23";
init_data(intToTimepoint(0))(22)(2, 1) <= x"1310";
init_data(intToTimepoint(1))(22)(2, 1) <= x"1310";
init_data(intToTimepoint(0))(23)(2, 1) <= x"0AFD";
init_data(intToTimepoint(1))(23)(2, 1) <= x"0AFD";
init_data(intToTimepoint(0))(24)(2, 1) <= x"2D93";
init_data(intToTimepoint(1))(24)(2, 1) <= x"2D93";
init_data(intToTimepoint(0))(25)(2, 1) <= x"278A";
init_data(intToTimepoint(1))(25)(2, 1) <= x"278A";
init_data(intToTimepoint(0))(26)(2, 1) <= x"2000";
init_data(intToTimepoint(1))(26)(2, 1) <= x"2000";
init_data(intToTimepoint(0))(27)(2, 1) <= x"17BD";
init_data(intToTimepoint(1))(27)(2, 1) <= x"17BD";
init_data(intToTimepoint(0))(28)(2, 1) <= x"0FA3";
init_data(intToTimepoint(1))(28)(2, 1) <= x"0FA3";
init_data(intToTimepoint(0))(29)(2, 1) <= x"0890";
init_data(intToTimepoint(1))(29)(2, 1) <= x"0890";
init_data(intToTimepoint(0))(30)(2, 1) <= x"2548";
init_data(intToTimepoint(1))(30)(2, 1) <= x"2548";
init_data(intToTimepoint(0))(31)(2, 1) <= x"2000";
init_data(intToTimepoint(1))(31)(2, 1) <= x"2000";
init_data(intToTimepoint(0))(32)(2, 1) <= x"1971";
init_data(intToTimepoint(1))(32)(2, 1) <= x"1971";
init_data(intToTimepoint(0))(33)(2, 1) <= x"1258";
init_data(intToTimepoint(1))(33)(2, 1) <= x"1258";
init_data(intToTimepoint(0))(34)(2, 1) <= x"0B84";
init_data(intToTimepoint(1))(34)(2, 1) <= x"0B84";
init_data(intToTimepoint(0))(35)(2, 1) <= x"05BF";
init_data(intToTimepoint(1))(35)(2, 1) <= x"05BF";
init_data(intToTimepoint(0))(0)(2, 2) <= x"0AFD";
init_data(intToTimepoint(1))(0)(2, 2) <= x"0AFD";
init_data(intToTimepoint(0))(1)(2, 2) <= x"0890";
init_data(intToTimepoint(1))(1)(2, 2) <= x"0890";
init_data(intToTimepoint(0))(2)(2, 2) <= x"05BF";
init_data(intToTimepoint(1))(2)(2, 2) <= x"05BF";
init_data(intToTimepoint(0))(3)(2, 2) <= x"0309";
init_data(intToTimepoint(1))(3)(2, 2) <= x"0309";
init_data(intToTimepoint(0))(4)(2, 2) <= x"00F5";
init_data(intToTimepoint(1))(4)(2, 2) <= x"00F5";
init_data(intToTimepoint(0))(5)(2, 2) <= x"0004";
init_data(intToTimepoint(1))(5)(2, 2) <= x"0004";
init_data(intToTimepoint(0))(6)(2, 2) <= x"1310";
init_data(intToTimepoint(1))(6)(2, 2) <= x"1310";
init_data(intToTimepoint(0))(7)(2, 2) <= x"0FA3";
init_data(intToTimepoint(1))(7)(2, 2) <= x"0FA3";
init_data(intToTimepoint(0))(8)(2, 2) <= x"0B84";
init_data(intToTimepoint(1))(8)(2, 2) <= x"0B84";
init_data(intToTimepoint(0))(9)(2, 2) <= x"0747";
init_data(intToTimepoint(1))(9)(2, 2) <= x"0747";
init_data(intToTimepoint(0))(10)(2, 2) <= x"038E";
init_data(intToTimepoint(1))(10)(2, 2) <= x"038E";
init_data(intToTimepoint(0))(11)(2, 2) <= x"00F5";
init_data(intToTimepoint(1))(11)(2, 2) <= x"00F5";
init_data(intToTimepoint(0))(12)(2, 2) <= x"1C23";
init_data(intToTimepoint(1))(12)(2, 2) <= x"1C23";
init_data(intToTimepoint(0))(13)(2, 2) <= x"17BD";
init_data(intToTimepoint(1))(13)(2, 2) <= x"17BD";
init_data(intToTimepoint(0))(14)(2, 2) <= x"1258";
init_data(intToTimepoint(1))(14)(2, 2) <= x"1258";
init_data(intToTimepoint(0))(15)(2, 2) <= x"0C9E";
init_data(intToTimepoint(1))(15)(2, 2) <= x"0C9E";
init_data(intToTimepoint(0))(16)(2, 2) <= x"0747";
init_data(intToTimepoint(1))(16)(2, 2) <= x"0747";
init_data(intToTimepoint(0))(17)(2, 2) <= x"0309";
init_data(intToTimepoint(1))(17)(2, 2) <= x"0309";
init_data(intToTimepoint(0))(18)(2, 2) <= x"2548";
init_data(intToTimepoint(1))(18)(2, 2) <= x"2548";
init_data(intToTimepoint(0))(19)(2, 2) <= x"2000";
init_data(intToTimepoint(1))(19)(2, 2) <= x"2000";
init_data(intToTimepoint(0))(20)(2, 2) <= x"1971";
init_data(intToTimepoint(1))(20)(2, 2) <= x"1971";
init_data(intToTimepoint(0))(21)(2, 2) <= x"1258";
init_data(intToTimepoint(1))(21)(2, 2) <= x"1258";
init_data(intToTimepoint(0))(22)(2, 2) <= x"0B84";
init_data(intToTimepoint(1))(22)(2, 2) <= x"0B84";
init_data(intToTimepoint(0))(23)(2, 2) <= x"05BF";
init_data(intToTimepoint(1))(23)(2, 2) <= x"05BF";
init_data(intToTimepoint(0))(24)(2, 2) <= x"2D93";
init_data(intToTimepoint(1))(24)(2, 2) <= x"2D93";
init_data(intToTimepoint(0))(25)(2, 2) <= x"278A";
init_data(intToTimepoint(1))(25)(2, 2) <= x"278A";
init_data(intToTimepoint(0))(26)(2, 2) <= x"2000";
init_data(intToTimepoint(1))(26)(2, 2) <= x"2000";
init_data(intToTimepoint(0))(27)(2, 2) <= x"17BD";
init_data(intToTimepoint(1))(27)(2, 2) <= x"17BD";
init_data(intToTimepoint(0))(28)(2, 2) <= x"0FA3";
init_data(intToTimepoint(1))(28)(2, 2) <= x"0FA3";
init_data(intToTimepoint(0))(29)(2, 2) <= x"0890";
init_data(intToTimepoint(1))(29)(2, 2) <= x"0890";
init_data(intToTimepoint(0))(30)(2, 2) <= x"342D";
init_data(intToTimepoint(1))(30)(2, 2) <= x"342D";
init_data(intToTimepoint(0))(31)(2, 2) <= x"2D93";
init_data(intToTimepoint(1))(31)(2, 2) <= x"2D93";
init_data(intToTimepoint(0))(32)(2, 2) <= x"2548";
init_data(intToTimepoint(1))(32)(2, 2) <= x"2548";
init_data(intToTimepoint(0))(33)(2, 2) <= x"1C23";
init_data(intToTimepoint(1))(33)(2, 2) <= x"1C23";
init_data(intToTimepoint(0))(34)(2, 2) <= x"1310";
init_data(intToTimepoint(1))(34)(2, 2) <= x"1310";
init_data(intToTimepoint(0))(35)(2, 2) <= x"0AFD";
init_data(intToTimepoint(1))(35)(2, 2) <= x"0AFD";
init_data(intToTimepoint(0))(0)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(0)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(1)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(1)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(2)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(2)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(3)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(3)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(4)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(4)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(5)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(5)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(6)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(6)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(7)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(7)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(8)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(8)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(9)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(9)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(10)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(10)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(11)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(11)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(12)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(12)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(13)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(13)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(14)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(14)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(15)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(15)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(16)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(16)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(17)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(17)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(18)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(18)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(19)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(19)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(20)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(20)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(21)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(21)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(22)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(22)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(23)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(23)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(24)(2, 3) <= x"00F5";
init_data(intToTimepoint(1))(24)(2, 3) <= x"00F5";
init_data(intToTimepoint(0))(25)(2, 3) <= x"006A";
init_data(intToTimepoint(1))(25)(2, 3) <= x"006A";
init_data(intToTimepoint(0))(26)(2, 3) <= x"0009";
init_data(intToTimepoint(1))(26)(2, 3) <= x"0009";
init_data(intToTimepoint(0))(27)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(27)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(28)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(28)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(29)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(29)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(30)(2, 3) <= x"04BC";
init_data(intToTimepoint(1))(30)(2, 3) <= x"04BC";
init_data(intToTimepoint(0))(31)(2, 3) <= x"034A";
init_data(intToTimepoint(1))(31)(2, 3) <= x"034A";
init_data(intToTimepoint(0))(32)(2, 3) <= x"01BE";
init_data(intToTimepoint(1))(32)(2, 3) <= x"01BE";
init_data(intToTimepoint(0))(33)(2, 3) <= x"0081";
init_data(intToTimepoint(1))(33)(2, 3) <= x"0081";
init_data(intToTimepoint(0))(34)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(34)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(35)(2, 3) <= x"0000";
init_data(intToTimepoint(1))(35)(2, 3) <= x"0000";
init_data(intToTimepoint(0))(0)(3, 0) <= x"0081";
init_data(intToTimepoint(1))(0)(3, 0) <= x"0081";
init_data(intToTimepoint(0))(1)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(1)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(2)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(2)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(3)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(3)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(4)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(4)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(5)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(5)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(6)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(6)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(7)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(7)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(8)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(8)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(9)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(9)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(10)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(10)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(11)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(11)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(12)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(12)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(13)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(13)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(14)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(14)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(15)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(15)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(16)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(16)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(17)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(17)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(18)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(18)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(19)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(19)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(20)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(20)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(21)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(21)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(22)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(22)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(23)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(23)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(24)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(24)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(25)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(25)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(26)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(26)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(27)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(27)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(28)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(28)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(29)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(29)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(30)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(30)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(31)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(31)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(32)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(32)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(33)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(33)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(34)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(34)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(35)(3, 0) <= x"0000";
init_data(intToTimepoint(1))(35)(3, 0) <= x"0000";
init_data(intToTimepoint(0))(0)(3, 1) <= x"05BF";
init_data(intToTimepoint(1))(0)(3, 1) <= x"05BF";
init_data(intToTimepoint(0))(1)(3, 1) <= x"0166";
init_data(intToTimepoint(1))(1)(3, 1) <= x"0166";
init_data(intToTimepoint(0))(2)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(2)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(3)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(3)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(4)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(4)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(5)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(5)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(6)(3, 1) <= x"061C";
init_data(intToTimepoint(1))(6)(3, 1) <= x"061C";
init_data(intToTimepoint(0))(7)(3, 1) <= x"0190";
init_data(intToTimepoint(1))(7)(3, 1) <= x"0190";
init_data(intToTimepoint(0))(8)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(8)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(9)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(9)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(10)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(10)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(11)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(11)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(12)(3, 1) <= x"05BF";
init_data(intToTimepoint(1))(12)(3, 1) <= x"05BF";
init_data(intToTimepoint(0))(13)(3, 1) <= x"0166";
init_data(intToTimepoint(1))(13)(3, 1) <= x"0166";
init_data(intToTimepoint(0))(14)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(14)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(15)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(15)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(16)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(16)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(17)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(17)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(18)(3, 1) <= x"04BC";
init_data(intToTimepoint(1))(18)(3, 1) <= x"04BC";
init_data(intToTimepoint(0))(19)(3, 1) <= x"00F5";
init_data(intToTimepoint(1))(19)(3, 1) <= x"00F5";
init_data(intToTimepoint(0))(20)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(20)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(21)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(21)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(22)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(22)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(23)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(23)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(24)(3, 1) <= x"034A";
init_data(intToTimepoint(1))(24)(3, 1) <= x"034A";
init_data(intToTimepoint(0))(25)(3, 1) <= x"006A";
init_data(intToTimepoint(1))(25)(3, 1) <= x"006A";
init_data(intToTimepoint(0))(26)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(26)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(27)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(27)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(28)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(28)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(29)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(29)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(30)(3, 1) <= x"01BE";
init_data(intToTimepoint(1))(30)(3, 1) <= x"01BE";
init_data(intToTimepoint(0))(31)(3, 1) <= x"0009";
init_data(intToTimepoint(1))(31)(3, 1) <= x"0009";
init_data(intToTimepoint(0))(32)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(32)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(33)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(33)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(34)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(34)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(35)(3, 1) <= x"0000";
init_data(intToTimepoint(1))(35)(3, 1) <= x"0000";
init_data(intToTimepoint(0))(0)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(0)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(1)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(1)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(2)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(2)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(3)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(3)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(4)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(4)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(5)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(5)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(6)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(6)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(7)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(7)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(8)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(8)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(9)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(9)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(10)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(10)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(11)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(11)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(12)(3, 2) <= x"0081";
init_data(intToTimepoint(1))(12)(3, 2) <= x"0081";
init_data(intToTimepoint(0))(13)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(13)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(14)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(14)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(15)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(15)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(16)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(16)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(17)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(17)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(18)(3, 2) <= x"01BE";
init_data(intToTimepoint(1))(18)(3, 2) <= x"01BE";
init_data(intToTimepoint(0))(19)(3, 2) <= x"0009";
init_data(intToTimepoint(1))(19)(3, 2) <= x"0009";
init_data(intToTimepoint(0))(20)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(20)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(21)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(21)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(22)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(22)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(23)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(23)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(24)(3, 2) <= x"034A";
init_data(intToTimepoint(1))(24)(3, 2) <= x"034A";
init_data(intToTimepoint(0))(25)(3, 2) <= x"006A";
init_data(intToTimepoint(1))(25)(3, 2) <= x"006A";
init_data(intToTimepoint(0))(26)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(26)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(27)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(27)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(28)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(28)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(29)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(29)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(30)(3, 2) <= x"04BC";
init_data(intToTimepoint(1))(30)(3, 2) <= x"04BC";
init_data(intToTimepoint(0))(31)(3, 2) <= x"00F5";
init_data(intToTimepoint(1))(31)(3, 2) <= x"00F5";
init_data(intToTimepoint(0))(32)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(32)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(33)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(33)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(34)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(34)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(35)(3, 2) <= x"0000";
init_data(intToTimepoint(1))(35)(3, 2) <= x"0000";
init_data(intToTimepoint(0))(0)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(0)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(1)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(1)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(2)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(2)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(3)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(3)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(4)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(4)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(5)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(5)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(6)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(6)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(7)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(7)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(8)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(8)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(9)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(9)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(10)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(10)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(11)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(11)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(12)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(12)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(13)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(13)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(14)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(14)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(15)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(15)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(16)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(16)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(17)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(17)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(18)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(18)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(19)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(19)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(20)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(20)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(21)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(21)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(22)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(22)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(23)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(23)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(24)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(24)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(25)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(25)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(26)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(26)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(27)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(27)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(28)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(28)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(29)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(29)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(30)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(30)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(31)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(31)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(32)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(32)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(33)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(33)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(34)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(34)(3, 3) <= x"0000";
init_data(intToTimepoint(0))(35)(3, 3) <= x"0000";
init_data(intToTimepoint(1))(35)(3, 3) <= x"0000";
end behavioral;
